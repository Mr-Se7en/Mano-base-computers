--==============================================================================
=========================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY AC_controller IS
   PORT ( d0                : IN  std_logic;
          d2                : IN  std_logic;
          d3                : IN  std_logic;
          logisimClockTree0 : IN  std_logic_vector( 4 DOWNTO 0 );
          t5                : IN  std_logic;
          L                 : OUT std_logic );
END ENTITY AC_controller;
